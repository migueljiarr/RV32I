





<!DOCTYPE html>
<html lang="en">
  <head>
    <meta charset="utf-8">



  <link crossorigin="anonymous" href="https://assets-cdn.github.com/assets/frameworks-81a59bf26d881d29286674f6deefe779c444382fff322085b50ba455460ccae5.css" integrity="sha256-gaWb8m2IHSkoZnT23u/necREOC//MiCFtQukVUYMyuU=" media="all" rel="stylesheet" />
  <link crossorigin="anonymous" href="https://assets-cdn.github.com/assets/github-87d822aa41a2e50fc4a176f81e161236c98e01a8a4e8258b55acdeab81d58d35.css" integrity="sha256-h9giqkGi5Q/EoXb4HhYSNsmOAaik6CWLVazeq4HVjTU=" media="all" rel="stylesheet" />
  
  
  
  

  <meta name="viewport" content="width=device-width">
  
  <title>riscv-tomthumb/constants.vhd at master · maikmerten/riscv-tomthumb</title>
  <link rel="search" type="application/opensearchdescription+xml" href="/opensearch.xml" title="GitHub">
  <link rel="fluid-icon" href="https://github.com/fluidicon.png" title="GitHub">
  <meta property="fb:app_id" content="1401488693436528">

    
    <meta content="https://avatars1.githubusercontent.com/u/2611432?v=3&amp;s=400" property="og:image" /><meta content="GitHub" property="og:site_name" /><meta content="object" property="og:type" /><meta content="maikmerten/riscv-tomthumb" property="og:title" /><meta content="https://github.com/maikmerten/riscv-tomthumb" property="og:url" /><meta content="riscv-tomthumb - A small RISC-V RV32I core written in VHDL, intended as testbed for my personal VHDL learning" property="og:description" />

  <link rel="assets" href="https://assets-cdn.github.com/">
  <link rel="web-socket" href="wss://live.github.com/_sockets/VjI6MTY5Mzc5Mzg1OjcyZTY3NDhmYTRhOWQ3NTBlMDk3MDI2Y2ZlMmQ4MWRiZGYyYmNjNTA5YjI4ZTI3OWQwNTA5YTE4OWZkM2U5MzE=--eaa7b99b93d826ecf0feb56754c09c7e2e558a20">
  <meta name="pjax-timeout" content="1000">
  <link rel="sudo-modal" href="/sessions/sudo_modal">
  <meta name="request-id" content="C6B7:502D:91FBC7:D6AF49:591C1B52" data-pjax-transient>
  

  <meta name="selected-link" value="repo_source" data-pjax-transient>

  <meta name="google-site-verification" content="KT5gs8h0wvaagLKAVWq8bbeNwnZZK1r1XQysX3xurLU">
<meta name="google-site-verification" content="ZzhVyEFwb7w3e0-uOTltm8Jsck2F5StVihD0exw2fsA">
    <meta name="google-analytics" content="UA-3769691-2">

<meta content="collector.githubapp.com" name="octolytics-host" /><meta content="github" name="octolytics-app-id" /><meta content="https://collector.githubapp.com/github-external/browser_event" name="octolytics-event-url" /><meta content="C6B7:502D:91FBC7:D6AF49:591C1B52" name="octolytics-dimension-request_id" /><meta content="27913866" name="octolytics-actor-id" /><meta content="Agonesc" name="octolytics-actor-login" /><meta content="f81f2a10f550495686a49c6e2fa491837acbac4f5a3b5a3d0c6f73515bc31558" name="octolytics-actor-hash" />
<meta content="/&lt;user-name&gt;/&lt;repo-name&gt;/blob/show" data-pjax-transient="true" name="analytics-location" />




  <meta class="js-ga-set" name="dimension1" content="Logged In">


  

      <meta name="hostname" content="github.com">
  <meta name="user-login" content="Agonesc">

      <meta name="expected-hostname" content="github.com">
    <meta name="js-proxy-site-detection-payload" content="NWUwNjBlZDViMmEzY2ZiMmZhMTAyNjc3OWZhZTY0YzE1NWUzNWJlZjA0OTdjYjljMjc5Yzg0OTg4ZWI3YzVjZHx7InJlbW90ZV9hZGRyZXNzIjoiODcuMjIxLjIuOTQiLCJyZXF1ZXN0X2lkIjoiQzZCNzo1MDJEOjkxRkJDNzpENkFGNDk6NTkxQzFCNTIiLCJ0aW1lc3RhbXAiOjE0OTUwMTQyMjYsImhvc3QiOiJnaXRodWIuY29tIn0=">


  <meta name="html-safe-nonce" content="ff64c46d0e579a5e532801141c62fd77627b9da2">

  <meta http-equiv="x-pjax-version" content="598266a6dd8e4f61e16b355161b735cd">
  

    
  <meta name="description" content="riscv-tomthumb - A small RISC-V RV32I core written in VHDL, intended as testbed for my personal VHDL learning">
  <meta name="go-import" content="github.com/maikmerten/riscv-tomthumb git https://github.com/maikmerten/riscv-tomthumb.git">

  <meta content="2611432" name="octolytics-dimension-user_id" /><meta content="maikmerten" name="octolytics-dimension-user_login" /><meta content="57315384" name="octolytics-dimension-repository_id" /><meta content="maikmerten/riscv-tomthumb" name="octolytics-dimension-repository_nwo" /><meta content="true" name="octolytics-dimension-repository_public" /><meta content="false" name="octolytics-dimension-repository_is_fork" /><meta content="57315384" name="octolytics-dimension-repository_network_root_id" /><meta content="maikmerten/riscv-tomthumb" name="octolytics-dimension-repository_network_root_nwo" />
  <link href="https://github.com/maikmerten/riscv-tomthumb/commits/master.atom" rel="alternate" title="Recent Commits to riscv-tomthumb:master" type="application/atom+xml">


    <link rel="canonical" href="https://github.com/maikmerten/riscv-tomthumb/blob/master/src/vhdl/cpu/constants.vhd" data-pjax-transient>


  <meta name="browser-stats-url" content="https://api.github.com/_private/browser/stats">

  <meta name="browser-errors-url" content="https://api.github.com/_private/browser/errors">

  <link rel="mask-icon" href="https://assets-cdn.github.com/pinned-octocat.svg" color="#000000">
  <link rel="icon" type="image/x-icon" href="https://assets-cdn.github.com/favicon.ico">

<meta name="theme-color" content="#1e2327">


  <meta name="u2f-support" content="true">

  </head>

  <body class="logged-in env-production page-blob">
    



  <div class="position-relative js-header-wrapper ">
    <a href="#start-of-content" tabindex="1" class="accessibility-aid js-skip-to-content">Skip to content</a>
    <div id="js-pjax-loader-bar" class="pjax-loader-bar"><div class="progress"></div></div>

    
    
    



        
<div class="header" role="banner">
  <div class="container clearfix">
    <a class="header-logo-invertocat" href="https://github.com/" data-hotkey="g d" aria-label="Homepage" data-ga-click="Header, go to dashboard, icon:logo">
  <svg aria-hidden="true" class="octicon octicon-mark-github" height="32" version="1.1" viewBox="0 0 16 16" width="32"><path fill-rule="evenodd" d="M8 0C3.58 0 0 3.58 0 8c0 3.54 2.29 6.53 5.47 7.59.4.07.55-.17.55-.38 0-.19-.01-.82-.01-1.49-2.01.37-2.53-.49-2.69-.94-.09-.23-.48-.94-.82-1.13-.28-.15-.68-.52-.01-.53.63-.01 1.08.58 1.23.82.72 1.21 1.87.87 2.33.66.07-.52.28-.87.51-1.07-1.78-.2-3.64-.89-3.64-3.95 0-.87.31-1.59.82-2.15-.08-.2-.36-1.02.08-2.12 0 0 .67-.21 2.2.82.64-.18 1.32-.27 2-.27.68 0 1.36.09 2 .27 1.53-1.04 2.2-.82 2.2-.82.44 1.1.16 1.92.08 2.12.51.56.82 1.27.82 2.15 0 3.07-1.87 3.75-3.65 3.95.29.25.54.73.54 1.48 0 1.07-.01 1.93-.01 2.2 0 .21.15.46.55.38A8.013 8.013 0 0 0 16 8c0-4.42-3.58-8-8-8z"/></svg>
</a>


        <div class="header-search scoped-search site-scoped-search js-site-search" role="search">
  <!-- '"` --><!-- </textarea></xmp> --></option></form><form accept-charset="UTF-8" action="/maikmerten/riscv-tomthumb/search" class="js-site-search-form" data-scoped-search-url="/maikmerten/riscv-tomthumb/search" data-unscoped-search-url="/search" method="get"><div style="margin:0;padding:0;display:inline"><input name="utf8" type="hidden" value="&#x2713;" /></div>
    <label class="form-control header-search-wrapper js-chromeless-input-container">
        <a href="/maikmerten/riscv-tomthumb/blob/master/src/vhdl/cpu/constants.vhd" class="header-search-scope no-underline">This repository</a>
      <input type="text"
        class="form-control header-search-input js-site-search-focus js-site-search-field is-clearable"
        data-hotkey="s"
        name="q"
        value=""
        placeholder="Search"
        aria-label="Search this repository"
        data-unscoped-placeholder="Search GitHub"
        data-scoped-placeholder="Search"
        autocapitalize="off">
        <input type="hidden" class="js-site-search-type-field" name="type" >
    </label>
</form></div>


      <ul class="header-nav float-left" role="navigation">
        <li class="header-nav-item">
          <a href="/pulls" aria-label="Pull requests you created" class="js-selected-navigation-item header-nav-link" data-ga-click="Header, click, Nav menu - item:pulls context:user" data-hotkey="g p" data-selected-links="/pulls /pulls/assigned /pulls/mentioned /pulls">
            Pull requests
</a>        </li>
        <li class="header-nav-item">
          <a href="/issues" aria-label="Issues you created" class="js-selected-navigation-item header-nav-link" data-ga-click="Header, click, Nav menu - item:issues context:user" data-hotkey="g i" data-selected-links="/issues /issues/assigned /issues/mentioned /issues">
            Issues
</a>        </li>
          <li class="header-nav-item">
            <a class="header-nav-link" href="https://gist.github.com/" data-ga-click="Header, go to gist, text:gist">Gist</a>
          </li>
      </ul>

    
<ul class="header-nav user-nav float-right" id="user-links">
  <li class="header-nav-item">
    

  </li>

  <li class="header-nav-item dropdown js-menu-container">
    <a class="header-nav-link tooltipped tooltipped-s js-menu-target" href="/new"
       aria-label="Create new…"
       data-ga-click="Header, create new, icon:add">
      <svg aria-hidden="true" class="octicon octicon-plus float-left" height="16" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M12 9H7v5H5V9H0V7h5V2h2v5h5z"/></svg>
      <span class="dropdown-caret"></span>
    </a>

    <div class="dropdown-menu-content js-menu-content">
      <ul class="dropdown-menu dropdown-menu-sw">
        
<a class="dropdown-item" href="/new" data-ga-click="Header, create new repository">
  New repository
</a>

  <a class="dropdown-item" href="/new/import" data-ga-click="Header, import a repository">
    Import repository
  </a>

<a class="dropdown-item" href="https://gist.github.com/" data-ga-click="Header, create new gist">
  New gist
</a>

  <a class="dropdown-item" href="/organizations/new" data-ga-click="Header, create new organization">
    New organization
  </a>



  <div class="dropdown-divider"></div>
  <div class="dropdown-header">
    <span title="maikmerten/riscv-tomthumb">This repository</span>
  </div>
    <a class="dropdown-item" href="/maikmerten/riscv-tomthumb/issues/new" data-ga-click="Header, create new issue">
      New issue
    </a>

      </ul>
    </div>
  </li>

  <li class="header-nav-item dropdown js-menu-container">
    <a class="header-nav-link name tooltipped tooltipped-sw js-menu-target" href="/Agonesc"
       aria-label="View profile and more"
       data-ga-click="Header, show menu, icon:avatar">
      <img alt="@Agonesc" class="avatar" src="https://avatars1.githubusercontent.com/u/27913866?v=3&amp;s=40" height="20" width="20">
      <span class="dropdown-caret"></span>
    </a>

    <div class="dropdown-menu-content js-menu-content">
      <div class="dropdown-menu dropdown-menu-sw">
        <div class="dropdown-header header-nav-current-user css-truncate">
          Signed in as <strong class="css-truncate-target">Agonesc</strong>
        </div>

        <div class="dropdown-divider"></div>

        <a class="dropdown-item" href="/Agonesc" data-ga-click="Header, go to profile, text:your profile">
          Your profile
        </a>
        <a class="dropdown-item" href="/Agonesc?tab=stars" data-ga-click="Header, go to starred repos, text:your stars">
          Your stars
        </a>
        <a class="dropdown-item" href="/explore" data-ga-click="Header, go to explore, text:explore">
          Explore
        </a>
          <a class="dropdown-item" href="/integrations" data-ga-click="Header, go to integrations, text:integrations">
            Integrations
          </a>
        <a class="dropdown-item" href="https://help.github.com" data-ga-click="Header, go to help, text:help">
          Help
        </a>

        <div class="dropdown-divider"></div>

        <a class="dropdown-item" href="/settings/profile" data-ga-click="Header, go to settings, icon:settings">
          Settings
        </a>

        <!-- '"` --><!-- </textarea></xmp> --></option></form><form accept-charset="UTF-8" action="/logout" class="logout-form" method="post"><div style="margin:0;padding:0;display:inline"><input name="utf8" type="hidden" value="&#x2713;" /><input name="authenticity_token" type="hidden" value="mKKNb5B/hhDXyml6oH18/7dj6jkKgfBFonkzfqg6BL4Ik6W5B5Nm380AvS9MbnKlgjjW5j969MBRYbMh/ygr6Q==" /></div>
          <button type="submit" class="dropdown-item dropdown-signout" data-ga-click="Header, sign out, icon:logout">
            Sign out
          </button>
</form>      </div>
    </div>
  </li>
</ul>


    <!-- '"` --><!-- </textarea></xmp> --></option></form><form accept-charset="UTF-8" action="/logout" class="sr-only right-0" method="post"><div style="margin:0;padding:0;display:inline"><input name="utf8" type="hidden" value="&#x2713;" /><input name="authenticity_token" type="hidden" value="KSLJVKvuOKTQq2v/JD2lepxceOj8sxUWRTGEYNy9Sai5E+GCPALYa8phv6rILqsgqQdEN8lIEZO2KQQ/i69m/w==" /></div>
      <button type="submit" class="dropdown-item dropdown-signout" data-ga-click="Header, sign out, icon:logout">
        Sign out
      </button>
</form>  </div>
</div>


      

  </div>

  <div id="start-of-content" class="accessibility-aid"></div>

    <div id="js-flash-container">
</div>



  <div role="main">
        <div itemscope itemtype="http://schema.org/SoftwareSourceCode">
    <div id="js-repo-pjax-container" data-pjax-container>
        



    <div class="pagehead repohead instapaper_ignore readability-menu experiment-repo-nav">
      <div class="container repohead-details-container">

        <ul class="pagehead-actions">
  <li>
        <!-- '"` --><!-- </textarea></xmp> --></option></form><form accept-charset="UTF-8" action="/notifications/subscribe" class="js-social-container" data-autosubmit="true" data-remote="true" method="post"><div style="margin:0;padding:0;display:inline"><input name="utf8" type="hidden" value="&#x2713;" /><input name="authenticity_token" type="hidden" value="B++b0O/x0cxPOA/OFYNktUzZ4Ga7WMSpXMjOGZH1t5SlUvwgYQxID0PKJwzDE/DxDFt86OkKAs15TNkl61XuKg==" /></div>      <input class="form-control" id="repository_id" name="repository_id" type="hidden" value="57315384" />

        <div class="select-menu js-menu-container js-select-menu">
          <a href="/maikmerten/riscv-tomthumb/subscription"
            class="btn btn-sm btn-with-count select-menu-button js-menu-target" role="button" tabindex="0" aria-haspopup="true"
            data-ga-click="Repository, click Watch settings, action:blob#show">
            <span class="js-select-button">
                <svg aria-hidden="true" class="octicon octicon-eye" height="16" version="1.1" viewBox="0 0 16 16" width="16"><path fill-rule="evenodd" d="M8.06 2C3 2 0 8 0 8s3 6 8.06 6C13 14 16 8 16 8s-3-6-7.94-6zM8 12c-2.2 0-4-1.78-4-4 0-2.2 1.8-4 4-4 2.22 0 4 1.8 4 4 0 2.22-1.78 4-4 4zm2-4c0 1.11-.89 2-2 2-1.11 0-2-.89-2-2 0-1.11.89-2 2-2 1.11 0 2 .89 2 2z"/></svg>
                Watch
            </span>
          </a>
            <a class="social-count js-social-count"
              href="/maikmerten/riscv-tomthumb/watchers"
              aria-label="1 user is watching this repository">
              1
            </a>

        <div class="select-menu-modal-holder">
          <div class="select-menu-modal subscription-menu-modal js-menu-content">
            <div class="select-menu-header js-navigation-enable" tabindex="-1">
              <svg aria-label="Close" class="octicon octicon-x js-menu-close" height="16" role="img" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M7.48 8l3.75 3.75-1.48 1.48L6 9.48l-3.75 3.75-1.48-1.48L4.52 8 .77 4.25l1.48-1.48L6 6.52l3.75-3.75 1.48 1.48z"/></svg>
              <span class="select-menu-title">Notifications</span>
            </div>

              <div class="select-menu-list js-navigation-container" role="menu">

                <div class="select-menu-item js-navigation-item selected" role="menuitem" tabindex="0">
                  <svg aria-hidden="true" class="octicon octicon-check select-menu-item-icon" height="16" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M12 5l-8 8-4-4 1.5-1.5L4 10l6.5-6.5z"/></svg>
                  <div class="select-menu-item-text">
                    <input checked="checked" id="do_included" name="do" type="radio" value="included" />
                    <span class="select-menu-item-heading">Not watching</span>
                    <span class="description">Be notified when participating or @mentioned.</span>
                    <span class="js-select-button-text hidden-select-button-text">
                      <svg aria-hidden="true" class="octicon octicon-eye" height="16" version="1.1" viewBox="0 0 16 16" width="16"><path fill-rule="evenodd" d="M8.06 2C3 2 0 8 0 8s3 6 8.06 6C13 14 16 8 16 8s-3-6-7.94-6zM8 12c-2.2 0-4-1.78-4-4 0-2.2 1.8-4 4-4 2.22 0 4 1.8 4 4 0 2.22-1.78 4-4 4zm2-4c0 1.11-.89 2-2 2-1.11 0-2-.89-2-2 0-1.11.89-2 2-2 1.11 0 2 .89 2 2z"/></svg>
                      Watch
                    </span>
                  </div>
                </div>

                <div class="select-menu-item js-navigation-item " role="menuitem" tabindex="0">
                  <svg aria-hidden="true" class="octicon octicon-check select-menu-item-icon" height="16" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M12 5l-8 8-4-4 1.5-1.5L4 10l6.5-6.5z"/></svg>
                  <div class="select-menu-item-text">
                    <input id="do_subscribed" name="do" type="radio" value="subscribed" />
                    <span class="select-menu-item-heading">Watching</span>
                    <span class="description">Be notified of all conversations.</span>
                    <span class="js-select-button-text hidden-select-button-text">
                      <svg aria-hidden="true" class="octicon octicon-eye" height="16" version="1.1" viewBox="0 0 16 16" width="16"><path fill-rule="evenodd" d="M8.06 2C3 2 0 8 0 8s3 6 8.06 6C13 14 16 8 16 8s-3-6-7.94-6zM8 12c-2.2 0-4-1.78-4-4 0-2.2 1.8-4 4-4 2.22 0 4 1.8 4 4 0 2.22-1.78 4-4 4zm2-4c0 1.11-.89 2-2 2-1.11 0-2-.89-2-2 0-1.11.89-2 2-2 1.11 0 2 .89 2 2z"/></svg>
                        Unwatch
                    </span>
                  </div>
                </div>

                <div class="select-menu-item js-navigation-item " role="menuitem" tabindex="0">
                  <svg aria-hidden="true" class="octicon octicon-check select-menu-item-icon" height="16" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M12 5l-8 8-4-4 1.5-1.5L4 10l6.5-6.5z"/></svg>
                  <div class="select-menu-item-text">
                    <input id="do_ignore" name="do" type="radio" value="ignore" />
                    <span class="select-menu-item-heading">Ignoring</span>
                    <span class="description">Never be notified.</span>
                    <span class="js-select-button-text hidden-select-button-text">
                      <svg aria-hidden="true" class="octicon octicon-mute" height="16" version="1.1" viewBox="0 0 16 16" width="16"><path fill-rule="evenodd" d="M8 2.81v10.38c0 .67-.81 1-1.28.53L3 10H1c-.55 0-1-.45-1-1V7c0-.55.45-1 1-1h2l3.72-3.72C7.19 1.81 8 2.14 8 2.81zm7.53 3.22l-1.06-1.06-1.97 1.97-1.97-1.97-1.06 1.06L11.44 8 9.47 9.97l1.06 1.06 1.97-1.97 1.97 1.97 1.06-1.06L13.56 8l1.97-1.97z"/></svg>
                        Stop ignoring
                    </span>
                  </div>
                </div>

              </div>

            </div>
          </div>
        </div>
</form>
  </li>

  <li>
      <div class="js-toggler-container js-social-container starring-container ">
    <!-- '"` --><!-- </textarea></xmp> --></option></form><form accept-charset="UTF-8" action="/maikmerten/riscv-tomthumb/unstar" class="starred" data-remote="true" method="post"><div style="margin:0;padding:0;display:inline"><input name="utf8" type="hidden" value="&#x2713;" /><input name="authenticity_token" type="hidden" value="ZSXqaryqj4VzABj2ZCh/irZAGzrzk9ZFxnwfyygTk4VwNwiGYq31v2AUQMTiw47J+4u9VleEVFCVZvWpO6PlTg==" /></div>
      <button
        type="submit"
        class="btn btn-sm btn-with-count js-toggler-target"
        aria-label="Unstar this repository" title="Unstar maikmerten/riscv-tomthumb"
        data-ga-click="Repository, click unstar button, action:blob#show; text:Unstar">
        <svg aria-hidden="true" class="octicon octicon-star" height="16" version="1.1" viewBox="0 0 14 16" width="14"><path fill-rule="evenodd" d="M14 6l-4.9-.64L7 1 4.9 5.36 0 6l3.6 3.26L2.67 14 7 11.67 11.33 14l-.93-4.74z"/></svg>
        Unstar
      </button>
        <a class="social-count js-social-count" href="/maikmerten/riscv-tomthumb/stargazers"
           aria-label="5 users starred this repository">
          5
        </a>
</form>
    <!-- '"` --><!-- </textarea></xmp> --></option></form><form accept-charset="UTF-8" action="/maikmerten/riscv-tomthumb/star" class="unstarred" data-remote="true" method="post"><div style="margin:0;padding:0;display:inline"><input name="utf8" type="hidden" value="&#x2713;" /><input name="authenticity_token" type="hidden" value="yypWtPB4XOBFTw1oClEwtP3JiqieU/tZHWQ22fCFe6paZcth+LSZCZZWVZIiqPP01uQ3efE6sGlNI0JFdnmKGA==" /></div>
      <button
        type="submit"
        class="btn btn-sm btn-with-count js-toggler-target"
        aria-label="Star this repository" title="Star maikmerten/riscv-tomthumb"
        data-ga-click="Repository, click star button, action:blob#show; text:Star">
        <svg aria-hidden="true" class="octicon octicon-star" height="16" version="1.1" viewBox="0 0 14 16" width="14"><path fill-rule="evenodd" d="M14 6l-4.9-.64L7 1 4.9 5.36 0 6l3.6 3.26L2.67 14 7 11.67 11.33 14l-.93-4.74z"/></svg>
        Star
      </button>
        <a class="social-count js-social-count" href="/maikmerten/riscv-tomthumb/stargazers"
           aria-label="5 users starred this repository">
          5
        </a>
</form>  </div>

  </li>

  <li>
          <!-- '"` --><!-- </textarea></xmp> --></option></form><form accept-charset="UTF-8" action="/maikmerten/riscv-tomthumb/fork" class="btn-with-count" method="post"><div style="margin:0;padding:0;display:inline"><input name="utf8" type="hidden" value="&#x2713;" /><input name="authenticity_token" type="hidden" value="pvZtVk3Nizkl3CqAam6ZI+enDFgbHfQnIxW2ES8zgTltLfdAco2zZwG3P8F1Fy1UWlNA2PMZ+LuM8clrXP2EtA==" /></div>
            <button
                type="submit"
                class="btn btn-sm btn-with-count"
                data-ga-click="Repository, show fork modal, action:blob#show; text:Fork"
                title="Fork your own copy of maikmerten/riscv-tomthumb to your account"
                aria-label="Fork your own copy of maikmerten/riscv-tomthumb to your account">
              <svg aria-hidden="true" class="octicon octicon-repo-forked" height="16" version="1.1" viewBox="0 0 10 16" width="10"><path fill-rule="evenodd" d="M8 1a1.993 1.993 0 0 0-1 3.72V6L5 8 3 6V4.72A1.993 1.993 0 0 0 2 1a1.993 1.993 0 0 0-1 3.72V6.5l3 3v1.78A1.993 1.993 0 0 0 5 15a1.993 1.993 0 0 0 1-3.72V9.5l3-3V4.72A1.993 1.993 0 0 0 8 1zM2 4.2C1.34 4.2.8 3.65.8 3c0-.65.55-1.2 1.2-1.2.65 0 1.2.55 1.2 1.2 0 .65-.55 1.2-1.2 1.2zm3 10c-.66 0-1.2-.55-1.2-1.2 0-.65.55-1.2 1.2-1.2.65 0 1.2.55 1.2 1.2 0 .65-.55 1.2-1.2 1.2zm3-10c-.66 0-1.2-.55-1.2-1.2 0-.65.55-1.2 1.2-1.2.65 0 1.2.55 1.2 1.2 0 .65-.55 1.2-1.2 1.2z"/></svg>
              Fork
            </button>
</form>
    <a href="/maikmerten/riscv-tomthumb/network" class="social-count"
       aria-label="1 user forked this repository">
      1
    </a>
  </li>
</ul>

        <h1 class="public ">
  <svg aria-hidden="true" class="octicon octicon-repo" height="16" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M4 9H3V8h1v1zm0-3H3v1h1V6zm0-2H3v1h1V4zm0-2H3v1h1V2zm8-1v12c0 .55-.45 1-1 1H6v2l-1.5-1.5L3 16v-2H1c-.55 0-1-.45-1-1V1c0-.55.45-1 1-1h10c.55 0 1 .45 1 1zm-1 10H1v2h2v-1h3v1h5v-2zm0-10H2v9h9V1z"/></svg>
  <span class="author" itemprop="author"><a href="/maikmerten" class="url fn" rel="author">maikmerten</a></span><!--
--><span class="path-divider">/</span><!--
--><strong itemprop="name"><a href="/maikmerten/riscv-tomthumb" data-pjax="#js-repo-pjax-container">riscv-tomthumb</a></strong>

</h1>

      </div>
      <div class="container">
        
<nav class="reponav js-repo-nav js-sidenav-container-pjax"
     itemscope
     itemtype="http://schema.org/BreadcrumbList"
     role="navigation"
     data-pjax="#js-repo-pjax-container">

  <span itemscope itemtype="http://schema.org/ListItem" itemprop="itemListElement">
    <a href="/maikmerten/riscv-tomthumb" class="js-selected-navigation-item selected reponav-item" data-hotkey="g c" data-selected-links="repo_source repo_downloads repo_commits repo_releases repo_tags repo_branches /maikmerten/riscv-tomthumb" itemprop="url">
      <svg aria-hidden="true" class="octicon octicon-code" height="16" version="1.1" viewBox="0 0 14 16" width="14"><path fill-rule="evenodd" d="M9.5 3L8 4.5 11.5 8 8 11.5 9.5 13 14 8 9.5 3zm-5 0L0 8l4.5 5L6 11.5 2.5 8 6 4.5 4.5 3z"/></svg>
      <span itemprop="name">Code</span>
      <meta itemprop="position" content="1">
</a>  </span>

    <span itemscope itemtype="http://schema.org/ListItem" itemprop="itemListElement">
      <a href="/maikmerten/riscv-tomthumb/issues" class="js-selected-navigation-item reponav-item" data-hotkey="g i" data-selected-links="repo_issues repo_labels repo_milestones /maikmerten/riscv-tomthumb/issues" itemprop="url">
        <svg aria-hidden="true" class="octicon octicon-issue-opened" height="16" version="1.1" viewBox="0 0 14 16" width="14"><path fill-rule="evenodd" d="M7 2.3c3.14 0 5.7 2.56 5.7 5.7s-2.56 5.7-5.7 5.7A5.71 5.71 0 0 1 1.3 8c0-3.14 2.56-5.7 5.7-5.7zM7 1C3.14 1 0 4.14 0 8s3.14 7 7 7 7-3.14 7-7-3.14-7-7-7zm1 3H6v5h2V4zm0 6H6v2h2v-2z"/></svg>
        <span itemprop="name">Issues</span>
        <span class="Counter">0</span>
        <meta itemprop="position" content="2">
</a>    </span>

  <span itemscope itemtype="http://schema.org/ListItem" itemprop="itemListElement">
    <a href="/maikmerten/riscv-tomthumb/pulls" class="js-selected-navigation-item reponav-item" data-hotkey="g p" data-selected-links="repo_pulls /maikmerten/riscv-tomthumb/pulls" itemprop="url">
      <svg aria-hidden="true" class="octicon octicon-git-pull-request" height="16" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M11 11.28V5c-.03-.78-.34-1.47-.94-2.06C9.46 2.35 8.78 2.03 8 2H7V0L4 3l3 3V4h1c.27.02.48.11.69.31.21.2.3.42.31.69v6.28A1.993 1.993 0 0 0 10 15a1.993 1.993 0 0 0 1-3.72zm-1 2.92c-.66 0-1.2-.55-1.2-1.2 0-.65.55-1.2 1.2-1.2.65 0 1.2.55 1.2 1.2 0 .65-.55 1.2-1.2 1.2zM4 3c0-1.11-.89-2-2-2a1.993 1.993 0 0 0-1 3.72v6.56A1.993 1.993 0 0 0 2 15a1.993 1.993 0 0 0 1-3.72V4.72c.59-.34 1-.98 1-1.72zm-.8 10c0 .66-.55 1.2-1.2 1.2-.65 0-1.2-.55-1.2-1.2 0-.65.55-1.2 1.2-1.2.65 0 1.2.55 1.2 1.2zM2 4.2C1.34 4.2.8 3.65.8 3c0-.65.55-1.2 1.2-1.2.65 0 1.2.55 1.2 1.2 0 .65-.55 1.2-1.2 1.2z"/></svg>
      <span itemprop="name">Pull requests</span>
      <span class="Counter">0</span>
      <meta itemprop="position" content="3">
</a>  </span>

    <a href="/maikmerten/riscv-tomthumb/projects" class="js-selected-navigation-item reponav-item" data-selected-links="repo_projects new_repo_project repo_project /maikmerten/riscv-tomthumb/projects">
      <svg aria-hidden="true" class="octicon octicon-project" height="16" version="1.1" viewBox="0 0 15 16" width="15"><path fill-rule="evenodd" d="M10 12h3V2h-3v10zm-4-2h3V2H6v8zm-4 4h3V2H2v12zm-1 1h13V1H1v14zM14 0H1a1 1 0 0 0-1 1v14a1 1 0 0 0 1 1h13a1 1 0 0 0 1-1V1a1 1 0 0 0-1-1z"/></svg>
      Projects
      <span class="Counter" >0</span>
</a>
    <a href="/maikmerten/riscv-tomthumb/wiki" class="js-selected-navigation-item reponav-item" data-hotkey="g w" data-selected-links="repo_wiki /maikmerten/riscv-tomthumb/wiki">
      <svg aria-hidden="true" class="octicon octicon-book" height="16" version="1.1" viewBox="0 0 16 16" width="16"><path fill-rule="evenodd" d="M3 5h4v1H3V5zm0 3h4V7H3v1zm0 2h4V9H3v1zm11-5h-4v1h4V5zm0 2h-4v1h4V7zm0 2h-4v1h4V9zm2-6v9c0 .55-.45 1-1 1H9.5l-1 1-1-1H2c-.55 0-1-.45-1-1V3c0-.55.45-1 1-1h5.5l1 1 1-1H15c.55 0 1 .45 1 1zm-8 .5L7.5 3H2v9h6V3.5zm7-.5H9.5l-.5.5V12h6V3z"/></svg>
      Wiki
</a>


  <a href="/maikmerten/riscv-tomthumb/pulse" class="js-selected-navigation-item reponav-item" data-selected-links="pulse /maikmerten/riscv-tomthumb/pulse">
    <svg aria-hidden="true" class="octicon octicon-pulse" height="16" version="1.1" viewBox="0 0 14 16" width="14"><path fill-rule="evenodd" d="M11.5 8L8.8 5.4 6.6 8.5 5.5 1.6 2.38 8H0v2h3.6l.9-1.8.9 5.4L9 8.5l1.6 1.5H14V8z"/></svg>
    Pulse
</a>
  <a href="/maikmerten/riscv-tomthumb/graphs" class="js-selected-navigation-item reponav-item" data-selected-links="repo_graphs repo_contributors /maikmerten/riscv-tomthumb/graphs">
    <svg aria-hidden="true" class="octicon octicon-graph" height="16" version="1.1" viewBox="0 0 16 16" width="16"><path fill-rule="evenodd" d="M16 14v1H0V0h1v14h15zM5 13H3V8h2v5zm4 0H7V3h2v10zm4 0h-2V6h2v7z"/></svg>
    Graphs
</a>

</nav>

      </div>
    </div>

<div class="container new-discussion-timeline experiment-repo-nav">
  <div class="repository-content">

    
          

<a href="/maikmerten/riscv-tomthumb/blob/af14d0552896e5ad6751808b6df34033ab534628/src/vhdl/cpu/constants.vhd" class="d-none js-permalink-shortcut" data-hotkey="y">Permalink</a>

<!-- blob contrib key: blob_contributors:v21:2b5cbf1f4f02eed7a207dd3f22449b0e -->

<div class="file-navigation js-zeroclipboard-container">
  
<div class="select-menu branch-select-menu js-menu-container js-select-menu float-left">
  <button class=" btn btn-sm select-menu-button js-menu-target css-truncate" data-hotkey="w"
    
    type="button" aria-label="Switch branches or tags" tabindex="0" aria-haspopup="true">
      <i>Branch:</i>
      <span class="js-select-button css-truncate-target">master</span>
  </button>

  <div class="select-menu-modal-holder js-menu-content js-navigation-container" data-pjax>

    <div class="select-menu-modal">
      <div class="select-menu-header">
        <svg aria-label="Close" class="octicon octicon-x js-menu-close" height="16" role="img" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M7.48 8l3.75 3.75-1.48 1.48L6 9.48l-3.75 3.75-1.48-1.48L4.52 8 .77 4.25l1.48-1.48L6 6.52l3.75-3.75 1.48 1.48z"/></svg>
        <span class="select-menu-title">Switch branches/tags</span>
      </div>

      <div class="select-menu-filters">
        <div class="select-menu-text-filter">
          <input type="text" aria-label="Filter branches/tags" id="context-commitish-filter-field" class="form-control js-filterable-field js-navigation-enable" placeholder="Filter branches/tags">
        </div>
        <div class="select-menu-tabs">
          <ul>
            <li class="select-menu-tab">
              <a href="#" data-tab-filter="branches" data-filter-placeholder="Filter branches/tags" class="js-select-menu-tab" role="tab">Branches</a>
            </li>
            <li class="select-menu-tab">
              <a href="#" data-tab-filter="tags" data-filter-placeholder="Find a tag…" class="js-select-menu-tab" role="tab">Tags</a>
            </li>
          </ul>
        </div>
      </div>

      <div class="select-menu-list select-menu-tab-bucket js-select-menu-tab-bucket" data-tab-filter="branches" role="menu">

        <div data-filterable-for="context-commitish-filter-field" data-filterable-type="substring">


            <a class="select-menu-item js-navigation-item js-navigation-open "
               href="/maikmerten/riscv-tomthumb/blob/alulight/src/vhdl/cpu/constants.vhd"
               data-name="alulight"
               data-skip-pjax="true"
               rel="nofollow">
              <svg aria-hidden="true" class="octicon octicon-check select-menu-item-icon" height="16" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M12 5l-8 8-4-4 1.5-1.5L4 10l6.5-6.5z"/></svg>
              <span class="select-menu-item-text css-truncate-target js-select-menu-filter-text">
                alulight
              </span>
            </a>
            <a class="select-menu-item js-navigation-item js-navigation-open "
               href="/maikmerten/riscv-tomthumb/blob/interrupts/src/vhdl/cpu/constants.vhd"
               data-name="interrupts"
               data-skip-pjax="true"
               rel="nofollow">
              <svg aria-hidden="true" class="octicon octicon-check select-menu-item-icon" height="16" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M12 5l-8 8-4-4 1.5-1.5L4 10l6.5-6.5z"/></svg>
              <span class="select-menu-item-text css-truncate-target js-select-menu-filter-text">
                interrupts
              </span>
            </a>
            <a class="select-menu-item js-navigation-item js-navigation-open selected"
               href="/maikmerten/riscv-tomthumb/blob/master/src/vhdl/cpu/constants.vhd"
               data-name="master"
               data-skip-pjax="true"
               rel="nofollow">
              <svg aria-hidden="true" class="octicon octicon-check select-menu-item-icon" height="16" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M12 5l-8 8-4-4 1.5-1.5L4 10l6.5-6.5z"/></svg>
              <span class="select-menu-item-text css-truncate-target js-select-menu-filter-text">
                master
              </span>
            </a>
            <a class="select-menu-item js-navigation-item js-navigation-open "
               href="/maikmerten/riscv-tomthumb/blob/trap/src/vhdl/cpu/constants.vhd"
               data-name="trap"
               data-skip-pjax="true"
               rel="nofollow">
              <svg aria-hidden="true" class="octicon octicon-check select-menu-item-icon" height="16" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M12 5l-8 8-4-4 1.5-1.5L4 10l6.5-6.5z"/></svg>
              <span class="select-menu-item-text css-truncate-target js-select-menu-filter-text">
                trap
              </span>
            </a>
        </div>

          <div class="select-menu-no-results">Nothing to show</div>
      </div>

      <div class="select-menu-list select-menu-tab-bucket js-select-menu-tab-bucket" data-tab-filter="tags">
        <div data-filterable-for="context-commitish-filter-field" data-filterable-type="substring">


        </div>

        <div class="select-menu-no-results">Nothing to show</div>
      </div>

    </div>
  </div>
</div>

  <div class="BtnGroup float-right">
    <a href="/maikmerten/riscv-tomthumb/find/master"
          class="js-pjax-capture-input btn btn-sm BtnGroup-item"
          data-pjax
          data-hotkey="t">
      Find file
    </a>
    <button aria-label="Copy file path to clipboard" class="js-zeroclipboard btn btn-sm BtnGroup-item tooltipped tooltipped-s" data-copied-hint="Copied!" type="button">Copy path</button>
  </div>
  <div class="breadcrumb js-zeroclipboard-target">
    <span class="repo-root js-repo-root"><span class="js-path-segment"><a href="/maikmerten/riscv-tomthumb"><span>riscv-tomthumb</span></a></span></span><span class="separator">/</span><span class="js-path-segment"><a href="/maikmerten/riscv-tomthumb/tree/master/src"><span>src</span></a></span><span class="separator">/</span><span class="js-path-segment"><a href="/maikmerten/riscv-tomthumb/tree/master/src/vhdl"><span>vhdl</span></a></span><span class="separator">/</span><span class="js-path-segment"><a href="/maikmerten/riscv-tomthumb/tree/master/src/vhdl/cpu"><span>cpu</span></a></span><span class="separator">/</span><strong class="final-path">constants.vhd</strong>
  </div>
</div>



  <div class="commit-tease">
      <span class="float-right">
        <a class="commit-tease-sha" href="/maikmerten/riscv-tomthumb/commit/3db0712c823eddefcd60a237cd6fda841cef44f3" data-pjax>
          3db0712
        </a>
        <relative-time datetime="2016-09-07T18:04:01Z">Sep 7, 2016</relative-time>
      </span>
      <div>
        <img alt="@maikmerten" class="avatar" height="20" src="https://avatars2.githubusercontent.com/u/2611432?v=3&amp;s=40" width="20" />
        <a href="/maikmerten" class="user-mention" rel="author">maikmerten</a>
          <a href="/maikmerten/riscv-tomthumb/commit/3db0712c823eddefcd60a237cd6fda841cef44f3" class="message" data-pjax="true" title="remove some unused PCU ops">remove some unused PCU ops</a>
      </div>

    <div class="commit-tease-contributors">
      <button type="button" class="btn-link muted-link contributors-toggle" data-facebox="#blob_contributors_box">
        <strong>1</strong>
         contributor
      </button>
      
    </div>

    <div id="blob_contributors_box" style="display:none">
      <h2 class="facebox-header" data-facebox-id="facebox-header">Users who have contributed to this file</h2>
      <ul class="facebox-user-list" data-facebox-id="facebox-description">
          <li class="facebox-user-list-item">
            <img alt="@maikmerten" height="24" src="https://avatars0.githubusercontent.com/u/2611432?v=3&amp;s=48" width="24" />
            <a href="/maikmerten">maikmerten</a>
          </li>
      </ul>
    </div>
  </div>

<div class="file">
  <div class="file-header">
  <div class="file-actions">

    <div class="BtnGroup">
      <a href="/maikmerten/riscv-tomthumb/raw/master/src/vhdl/cpu/constants.vhd" class="btn btn-sm BtnGroup-item" id="raw-url">Raw</a>
        <a href="/maikmerten/riscv-tomthumb/blame/master/src/vhdl/cpu/constants.vhd" class="btn btn-sm js-update-url-with-hash BtnGroup-item" data-hotkey="b">Blame</a>
      <a href="/maikmerten/riscv-tomthumb/commits/master/src/vhdl/cpu/constants.vhd" class="btn btn-sm BtnGroup-item" rel="nofollow">History</a>
    </div>

        <a class="btn-octicon tooltipped tooltipped-nw"
           href="https://desktop.github.com"
           aria-label="Open this file in GitHub Desktop"
           data-ga-click="Repository, open with desktop, type:windows">
            <svg aria-hidden="true" class="octicon octicon-device-desktop" height="16" version="1.1" viewBox="0 0 16 16" width="16"><path fill-rule="evenodd" d="M15 2H1c-.55 0-1 .45-1 1v9c0 .55.45 1 1 1h5.34c-.25.61-.86 1.39-2.34 2h8c-1.48-.61-2.09-1.39-2.34-2H15c.55 0 1-.45 1-1V3c0-.55-.45-1-1-1zm0 9H1V3h14v8z"/></svg>
        </a>

        <!-- '"` --><!-- </textarea></xmp> --></option></form><form accept-charset="UTF-8" action="/maikmerten/riscv-tomthumb/edit/master/src/vhdl/cpu/constants.vhd" class="inline-form js-update-url-with-hash" method="post"><div style="margin:0;padding:0;display:inline"><input name="utf8" type="hidden" value="&#x2713;" /><input name="authenticity_token" type="hidden" value="ZXQJhSQVxjzQtyNL4SrPa8RmZr32/S3H4WMZSupptcg3fK6OThCJGsu7vdYdB8onRJ+aymqwF9Jd/KQQwM5Z9Q==" /></div>
          <button class="btn-octicon tooltipped tooltipped-nw" type="submit"
            aria-label="Fork this project and edit the file" data-hotkey="e" data-disable-with>
            <svg aria-hidden="true" class="octicon octicon-pencil" height="16" version="1.1" viewBox="0 0 14 16" width="14"><path fill-rule="evenodd" d="M0 12v3h3l8-8-3-3-8 8zm3 2H1v-2h1v1h1v1zm10.3-9.3L12 6 9 3l1.3-1.3a.996.996 0 0 1 1.41 0l1.59 1.59c.39.39.39 1.02 0 1.41z"/></svg>
          </button>
</form>        <!-- '"` --><!-- </textarea></xmp> --></option></form><form accept-charset="UTF-8" action="/maikmerten/riscv-tomthumb/delete/master/src/vhdl/cpu/constants.vhd" class="inline-form" method="post"><div style="margin:0;padding:0;display:inline"><input name="utf8" type="hidden" value="&#x2713;" /><input name="authenticity_token" type="hidden" value="fBVy7EvnQD8SMSL6KNadw646sOydS8mkRGGxeMBXOEsxCm1BkQD4JAlyIz3fOzlEAPg+31u/trpel5FKkWkbJg==" /></div>
          <button class="btn-octicon btn-octicon-danger tooltipped tooltipped-nw" type="submit"
            aria-label="Fork this project and delete the file" data-disable-with>
            <svg aria-hidden="true" class="octicon octicon-trashcan" height="16" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M11 2H9c0-.55-.45-1-1-1H5c-.55 0-1 .45-1 1H2c-.55 0-1 .45-1 1v1c0 .55.45 1 1 1v9c0 .55.45 1 1 1h7c.55 0 1-.45 1-1V5c.55 0 1-.45 1-1V3c0-.55-.45-1-1-1zm-1 12H3V5h1v8h1V5h1v8h1V5h1v8h1V5h1v9zm1-10H2V3h9v1z"/></svg>
          </button>
</form>  </div>

  <div class="file-info">
      158 lines (122 sloc)
      <span class="file-info-divider"></span>
    6.56 KB
  </div>
</div>

  

  <div itemprop="text" class="blob-wrapper data type-vhdl">
      <table class="highlight tab-size js-file-line-container" data-tab-size="8">
      <tr>
        <td id="L1" class="blob-num js-line-number" data-line-number="1"></td>
        <td id="LC1" class="blob-code blob-code-inner js-file-line"><span class="pl-k">library</span> IEEE;</td>
      </tr>
      <tr>
        <td id="L2" class="blob-num js-line-number" data-line-number="2"></td>
        <td id="LC2" class="blob-code blob-code-inner js-file-line"><span class="pl-k">use</span> IEEE.STD_LOGIC_1164.<span class="pl-k">all</span>;</td>
      </tr>
      <tr>
        <td id="L3" class="blob-num js-line-number" data-line-number="3"></td>
        <td id="LC3" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L4" class="blob-num js-line-number" data-line-number="4"></td>
        <td id="LC4" class="blob-code blob-code-inner js-file-line"><span class="pl-k">package</span> <span class="pl-en">constants</span> <span class="pl-k">is</span></td>
      </tr>
      <tr>
        <td id="L5" class="blob-num js-line-number" data-line-number="5"></td>
        <td id="LC5" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L6" class="blob-num js-line-number" data-line-number="6"></td>
        <td id="LC6" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> XLEN:	<span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">32</span>;</td>
      </tr>
      <tr>
        <td id="L7" class="blob-num js-line-number" data-line-number="7"></td>
        <td id="LC7" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> XLEN_ZERO: <span class="pl-c1">std_logic_vector</span>(XLEN<span class="pl-k">-</span><span class="pl-c1">1</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">X&quot;00000000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L8" class="blob-num js-line-number" data-line-number="8"></td>
        <td id="LC8" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> XLEN_ONE: <span class="pl-c1">std_logic_vector</span>(XLEN<span class="pl-k">-</span><span class="pl-c1">1</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">X&quot;00000001&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L9" class="blob-num js-line-number" data-line-number="9"></td>
        <td id="LC9" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L10" class="blob-num js-line-number" data-line-number="10"></td>
        <td id="LC10" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> RESET_VECTOR: 		<span class="pl-c1">std_logic_vector</span>(XLEN<span class="pl-k">-</span><span class="pl-c1">1</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">X&quot;00000000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L11" class="blob-num js-line-number" data-line-number="11"></td>
        <td id="LC11" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> TRAP_VECTOR:		<span class="pl-c1">std_logic_vector</span>(XLEN<span class="pl-k">-</span><span class="pl-c1">1</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">X&quot;00000004&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L12" class="blob-num js-line-number" data-line-number="12"></td>
        <td id="LC12" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> INTERRUPT_VECTOR:	<span class="pl-c1">std_logic_vector</span>(XLEN<span class="pl-k">-</span><span class="pl-c1">1</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">X&quot;00000008&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L13" class="blob-num js-line-number" data-line-number="13"></td>
        <td id="LC13" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L14" class="blob-num js-line-number" data-line-number="14"></td>
        <td id="LC14" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L15" class="blob-num js-line-number" data-line-number="15"></td>
        <td id="LC15" class="blob-code blob-code-inner js-file-line"><span class="pl-c"><span class="pl-c">--</span> Opcodes</span></td>
      </tr>
      <tr>
        <td id="L16" class="blob-num js-line-number" data-line-number="16"></td>
        <td id="LC16" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> OP_OP: 		<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;01100&quot;</span>; <span class="pl-c"><span class="pl-c">--</span> R-type</span></td>
      </tr>
      <tr>
        <td id="L17" class="blob-num js-line-number" data-line-number="17"></td>
        <td id="LC17" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> OP_CUSTOM0:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;00010&quot;</span>; <span class="pl-c"><span class="pl-c">--</span> R-type</span></td>
      </tr>
      <tr>
        <td id="L18" class="blob-num js-line-number" data-line-number="18"></td>
        <td id="LC18" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L19" class="blob-num js-line-number" data-line-number="19"></td>
        <td id="LC19" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> OP_JALR:		<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;11001&quot;</span>; <span class="pl-c"><span class="pl-c">--</span> I-type</span></td>
      </tr>
      <tr>
        <td id="L20" class="blob-num js-line-number" data-line-number="20"></td>
        <td id="LC20" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> OP_LOAD: 	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;00000&quot;</span>; <span class="pl-c"><span class="pl-c">--</span> I-type</span></td>
      </tr>
      <tr>
        <td id="L21" class="blob-num js-line-number" data-line-number="21"></td>
        <td id="LC21" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> OP_OPIMM: 	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;00100&quot;</span>; <span class="pl-c"><span class="pl-c">--</span> I-type</span></td>
      </tr>
      <tr>
        <td id="L22" class="blob-num js-line-number" data-line-number="22"></td>
        <td id="LC22" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> OP_SYSTEM: 	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;11100&quot;</span>; <span class="pl-c"><span class="pl-c">--</span> I-type</span></td>
      </tr>
      <tr>
        <td id="L23" class="blob-num js-line-number" data-line-number="23"></td>
        <td id="LC23" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> OP_MISCMEM: <span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;00011&quot;</span>; <span class="pl-c"><span class="pl-c">--</span> I-type?</span></td>
      </tr>
      <tr>
        <td id="L24" class="blob-num js-line-number" data-line-number="24"></td>
        <td id="LC24" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L25" class="blob-num js-line-number" data-line-number="25"></td>
        <td id="LC25" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> OP_STORE: 	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;01000&quot;</span>; <span class="pl-c"><span class="pl-c">--</span> S-type</span></td>
      </tr>
      <tr>
        <td id="L26" class="blob-num js-line-number" data-line-number="26"></td>
        <td id="LC26" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L27" class="blob-num js-line-number" data-line-number="27"></td>
        <td id="LC27" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> OP_BRANCH: 	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;11000&quot;</span>; <span class="pl-c"><span class="pl-c">--</span> SB-type</span></td>
      </tr>
      <tr>
        <td id="L28" class="blob-num js-line-number" data-line-number="28"></td>
        <td id="LC28" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L29" class="blob-num js-line-number" data-line-number="29"></td>
        <td id="LC29" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> OP_LUI: 		<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;01101&quot;</span>; <span class="pl-c"><span class="pl-c">--</span> U-type</span></td>
      </tr>
      <tr>
        <td id="L30" class="blob-num js-line-number" data-line-number="30"></td>
        <td id="LC30" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> OP_AUIPC: 	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;00101&quot;</span>; <span class="pl-c"><span class="pl-c">--</span> U-type</span></td>
      </tr>
      <tr>
        <td id="L31" class="blob-num js-line-number" data-line-number="31"></td>
        <td id="LC31" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L32" class="blob-num js-line-number" data-line-number="32"></td>
        <td id="LC32" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> OP_JAL: 		<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;11011&quot;</span>; <span class="pl-c"><span class="pl-c">--</span> UJ-type</span></td>
      </tr>
      <tr>
        <td id="L33" class="blob-num js-line-number" data-line-number="33"></td>
        <td id="LC33" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L34" class="blob-num js-line-number" data-line-number="34"></td>
        <td id="LC34" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_JALR:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L35" class="blob-num js-line-number" data-line-number="35"></td>
        <td id="LC35" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L36" class="blob-num js-line-number" data-line-number="36"></td>
        <td id="LC36" class="blob-code blob-code-inner js-file-line"><span class="pl-c"><span class="pl-c">--</span> Functions</span></td>
      </tr>
      <tr>
        <td id="L37" class="blob-num js-line-number" data-line-number="37"></td>
        <td id="LC37" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L38" class="blob-num js-line-number" data-line-number="38"></td>
        <td id="LC38" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_BEQ:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L39" class="blob-num js-line-number" data-line-number="39"></td>
        <td id="LC39" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_BNE:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;001&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L40" class="blob-num js-line-number" data-line-number="40"></td>
        <td id="LC40" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_BLT:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;100&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L41" class="blob-num js-line-number" data-line-number="41"></td>
        <td id="LC41" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_BGE:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;101&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L42" class="blob-num js-line-number" data-line-number="42"></td>
        <td id="LC42" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_BLTU:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;110&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L43" class="blob-num js-line-number" data-line-number="43"></td>
        <td id="LC43" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_BGEU:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;111&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L44" class="blob-num js-line-number" data-line-number="44"></td>
        <td id="LC44" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L45" class="blob-num js-line-number" data-line-number="45"></td>
        <td id="LC45" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_LB:		<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L46" class="blob-num js-line-number" data-line-number="46"></td>
        <td id="LC46" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_LH:		<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;001&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L47" class="blob-num js-line-number" data-line-number="47"></td>
        <td id="LC47" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_LW:		<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;010&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L48" class="blob-num js-line-number" data-line-number="48"></td>
        <td id="LC48" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_LBU:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;100&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L49" class="blob-num js-line-number" data-line-number="49"></td>
        <td id="LC49" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_LHU:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;101&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L50" class="blob-num js-line-number" data-line-number="50"></td>
        <td id="LC50" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L51" class="blob-num js-line-number" data-line-number="51"></td>
        <td id="LC51" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_SB:		<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L52" class="blob-num js-line-number" data-line-number="52"></td>
        <td id="LC52" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_SH:		<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;001&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L53" class="blob-num js-line-number" data-line-number="53"></td>
        <td id="LC53" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_SW:		<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;010&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L54" class="blob-num js-line-number" data-line-number="54"></td>
        <td id="LC54" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L55" class="blob-num js-line-number" data-line-number="55"></td>
        <td id="LC55" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_ADDI:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L56" class="blob-num js-line-number" data-line-number="56"></td>
        <td id="LC56" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_SLLI:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;001&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L57" class="blob-num js-line-number" data-line-number="57"></td>
        <td id="LC57" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_SLTI:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;010&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L58" class="blob-num js-line-number" data-line-number="58"></td>
        <td id="LC58" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_SLTIU:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;011&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L59" class="blob-num js-line-number" data-line-number="59"></td>
        <td id="LC59" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_XORI:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;100&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L60" class="blob-num js-line-number" data-line-number="60"></td>
        <td id="LC60" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_SRLI_SRAI:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;101&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L61" class="blob-num js-line-number" data-line-number="61"></td>
        <td id="LC61" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_ORI:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;110&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L62" class="blob-num js-line-number" data-line-number="62"></td>
        <td id="LC62" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_ANDI:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;111&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L63" class="blob-num js-line-number" data-line-number="63"></td>
        <td id="LC63" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L64" class="blob-num js-line-number" data-line-number="64"></td>
        <td id="LC64" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_ADD_SUB:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L65" class="blob-num js-line-number" data-line-number="65"></td>
        <td id="LC65" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_SLL:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;001&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L66" class="blob-num js-line-number" data-line-number="66"></td>
        <td id="LC66" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_SLT:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;010&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L67" class="blob-num js-line-number" data-line-number="67"></td>
        <td id="LC67" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_SLTU:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;011&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L68" class="blob-num js-line-number" data-line-number="68"></td>
        <td id="LC68" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_XOR:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;100&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L69" class="blob-num js-line-number" data-line-number="69"></td>
        <td id="LC69" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_SRL_SRA:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;101&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L70" class="blob-num js-line-number" data-line-number="70"></td>
        <td id="LC70" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_OR:		<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;110&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L71" class="blob-num js-line-number" data-line-number="71"></td>
        <td id="LC71" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_AND:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;111&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L72" class="blob-num js-line-number" data-line-number="72"></td>
        <td id="LC72" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L73" class="blob-num js-line-number" data-line-number="73"></td>
        <td id="LC73" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_FENCE:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L74" class="blob-num js-line-number" data-line-number="74"></td>
        <td id="LC74" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_FENCEI:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;001&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L75" class="blob-num js-line-number" data-line-number="75"></td>
        <td id="LC75" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L76" class="blob-num js-line-number" data-line-number="76"></td>
        <td id="LC76" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_SCALL_SBREAK:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L77" class="blob-num js-line-number" data-line-number="77"></td>
        <td id="LC77" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> FUNC_RD:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">2</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;010&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L78" class="blob-num js-line-number" data-line-number="78"></td>
        <td id="LC78" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L79" class="blob-num js-line-number" data-line-number="79"></td>
        <td id="LC79" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L80" class="blob-num js-line-number" data-line-number="80"></td>
        <td id="LC80" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R0:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;00000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L81" class="blob-num js-line-number" data-line-number="81"></td>
        <td id="LC81" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R1:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;00001&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L82" class="blob-num js-line-number" data-line-number="82"></td>
        <td id="LC82" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R2:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;00010&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L83" class="blob-num js-line-number" data-line-number="83"></td>
        <td id="LC83" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R3:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;00011&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L84" class="blob-num js-line-number" data-line-number="84"></td>
        <td id="LC84" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R4:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;00100&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L85" class="blob-num js-line-number" data-line-number="85"></td>
        <td id="LC85" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R5, T0:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;00101&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L86" class="blob-num js-line-number" data-line-number="86"></td>
        <td id="LC86" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R6, T1:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;00110&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L87" class="blob-num js-line-number" data-line-number="87"></td>
        <td id="LC87" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R7, T2:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;00111&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L88" class="blob-num js-line-number" data-line-number="88"></td>
        <td id="LC88" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R8:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;01000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L89" class="blob-num js-line-number" data-line-number="89"></td>
        <td id="LC89" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R9:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;01001&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L90" class="blob-num js-line-number" data-line-number="90"></td>
        <td id="LC90" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R10:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;01010&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L91" class="blob-num js-line-number" data-line-number="91"></td>
        <td id="LC91" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R11:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;01011&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L92" class="blob-num js-line-number" data-line-number="92"></td>
        <td id="LC92" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R12:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;01100&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L93" class="blob-num js-line-number" data-line-number="93"></td>
        <td id="LC93" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R13:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;01101&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L94" class="blob-num js-line-number" data-line-number="94"></td>
        <td id="LC94" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R14:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;01110&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L95" class="blob-num js-line-number" data-line-number="95"></td>
        <td id="LC95" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R15:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;01111&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L96" class="blob-num js-line-number" data-line-number="96"></td>
        <td id="LC96" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R16:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;10000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L97" class="blob-num js-line-number" data-line-number="97"></td>
        <td id="LC97" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R17:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;10001&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L98" class="blob-num js-line-number" data-line-number="98"></td>
        <td id="LC98" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R18:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;10010&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L99" class="blob-num js-line-number" data-line-number="99"></td>
        <td id="LC99" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R19:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;10011&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L100" class="blob-num js-line-number" data-line-number="100"></td>
        <td id="LC100" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R20:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;10100&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L101" class="blob-num js-line-number" data-line-number="101"></td>
        <td id="LC101" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R21:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;10101&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L102" class="blob-num js-line-number" data-line-number="102"></td>
        <td id="LC102" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R22:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;10110&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L103" class="blob-num js-line-number" data-line-number="103"></td>
        <td id="LC103" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R23:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;10111&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L104" class="blob-num js-line-number" data-line-number="104"></td>
        <td id="LC104" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R24:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;11000&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L105" class="blob-num js-line-number" data-line-number="105"></td>
        <td id="LC105" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R25:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;11001&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L106" class="blob-num js-line-number" data-line-number="106"></td>
        <td id="LC106" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R26:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;11010&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L107" class="blob-num js-line-number" data-line-number="107"></td>
        <td id="LC107" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R27:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;11011&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L108" class="blob-num js-line-number" data-line-number="108"></td>
        <td id="LC108" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R28:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;11100&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L109" class="blob-num js-line-number" data-line-number="109"></td>
        <td id="LC109" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R29:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;11101&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L110" class="blob-num js-line-number" data-line-number="110"></td>
        <td id="LC110" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R30:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;11110&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L111" class="blob-num js-line-number" data-line-number="111"></td>
        <td id="LC111" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> R31:	<span class="pl-c1">std_logic_vector</span>(<span class="pl-c1">4</span> <span class="pl-k">downto</span> <span class="pl-c1">0</span>) <span class="pl-k">:=</span> <span class="pl-c1">&quot;11111&quot;</span>;</td>
      </tr>
      <tr>
        <td id="L112" class="blob-num js-line-number" data-line-number="112"></td>
        <td id="LC112" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L113" class="blob-num js-line-number" data-line-number="113"></td>
        <td id="LC113" class="blob-code blob-code-inner js-file-line"><span class="pl-c"><span class="pl-c">--</span> muxer ports</span></td>
      </tr>
      <tr>
        <td id="L114" class="blob-num js-line-number" data-line-number="114"></td>
        <td id="LC114" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L115" class="blob-num js-line-number" data-line-number="115"></td>
        <td id="LC115" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_BUS_ADDR_PORTS: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">2</span>;</td>
      </tr>
      <tr>
        <td id="L116" class="blob-num js-line-number" data-line-number="116"></td>
        <td id="LC116" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_BUS_ADDR_PORT_ALU: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">0</span>;</td>
      </tr>
      <tr>
        <td id="L117" class="blob-num js-line-number" data-line-number="117"></td>
        <td id="LC117" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_BUS_ADDR_PORT_PC: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">1</span>;</td>
      </tr>
      <tr>
        <td id="L118" class="blob-num js-line-number" data-line-number="118"></td>
        <td id="LC118" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L119" class="blob-num js-line-number" data-line-number="119"></td>
        <td id="LC119" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_REG_DATA_PORTS: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">4</span>;</td>
      </tr>
      <tr>
        <td id="L120" class="blob-num js-line-number" data-line-number="120"></td>
        <td id="LC120" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_REG_DATA_PORT_ALU: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">0</span>;</td>
      </tr>
      <tr>
        <td id="L121" class="blob-num js-line-number" data-line-number="121"></td>
        <td id="LC121" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_REG_DATA_PORT_BUS: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">1</span>;</td>
      </tr>
      <tr>
        <td id="L122" class="blob-num js-line-number" data-line-number="122"></td>
        <td id="LC122" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_REG_DATA_PORT_IMM: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">2</span>;</td>
      </tr>
      <tr>
        <td id="L123" class="blob-num js-line-number" data-line-number="123"></td>
        <td id="LC123" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_REG_DATA_PORT_TRAPRET: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">3</span>;</td>
      </tr>
      <tr>
        <td id="L124" class="blob-num js-line-number" data-line-number="124"></td>
        <td id="LC124" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L125" class="blob-num js-line-number" data-line-number="125"></td>
        <td id="LC125" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_ALU_DAT1_PORTS: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">2</span>;</td>
      </tr>
      <tr>
        <td id="L126" class="blob-num js-line-number" data-line-number="126"></td>
        <td id="LC126" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_ALU_DAT1_PORT_S1: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">0</span>;</td>
      </tr>
      <tr>
        <td id="L127" class="blob-num js-line-number" data-line-number="127"></td>
        <td id="LC127" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_ALU_DAT1_PORT_PC: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">1</span>;</td>
      </tr>
      <tr>
        <td id="L128" class="blob-num js-line-number" data-line-number="128"></td>
        <td id="LC128" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L129" class="blob-num js-line-number" data-line-number="129"></td>
        <td id="LC129" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_ALU_DAT2_PORTS: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">3</span>;</td>
      </tr>
      <tr>
        <td id="L130" class="blob-num js-line-number" data-line-number="130"></td>
        <td id="LC130" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_ALU_DAT2_PORT_S2: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">0</span>;</td>
      </tr>
      <tr>
        <td id="L131" class="blob-num js-line-number" data-line-number="131"></td>
        <td id="LC131" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_ALU_DAT2_PORT_IMM: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">1</span>;</td>
      </tr>
      <tr>
        <td id="L132" class="blob-num js-line-number" data-line-number="132"></td>
        <td id="LC132" class="blob-code blob-code-inner js-file-line"><span class="pl-k">constant</span> MUX_ALU_DAT2_PORT_INSTLEN: <span class="pl-c1">integer</span> <span class="pl-k">:=</span> <span class="pl-c1">2</span>;</td>
      </tr>
      <tr>
        <td id="L133" class="blob-num js-line-number" data-line-number="133"></td>
        <td id="LC133" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L134" class="blob-num js-line-number" data-line-number="134"></td>
        <td id="LC134" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L135" class="blob-num js-line-number" data-line-number="135"></td>
        <td id="LC135" class="blob-code blob-code-inner js-file-line"><span class="pl-k">attribute</span> enum_encoding : <span class="pl-c1">string</span>;</td>
      </tr>
      <tr>
        <td id="L136" class="blob-num js-line-number" data-line-number="136"></td>
        <td id="LC136" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L137" class="blob-num js-line-number" data-line-number="137"></td>
        <td id="LC137" class="blob-code blob-code-inner js-file-line"><span class="pl-c"><span class="pl-c">--</span> ALU operations, signalled by decode unit</span></td>
      </tr>
      <tr>
        <td id="L138" class="blob-num js-line-number" data-line-number="138"></td>
        <td id="LC138" class="blob-code blob-code-inner js-file-line"><span class="pl-k">type</span> <span class="pl-en">aluops_t</span> <span class="pl-k">is</span> (ALU_ADD, ALU_SUB, ALU_AND, ALU_OR, ALU_XOR, ALU_SLT, ALU_SLTU, ALU_SLL, ALU_SRL, ALU_SRA);</td>
      </tr>
      <tr>
        <td id="L139" class="blob-num js-line-number" data-line-number="139"></td>
        <td id="LC139" class="blob-code blob-code-inner js-file-line"><span class="pl-c"><span class="pl-c">--</span>attribute enum_encoding of aluops_t : type is &quot;sequential&quot;;</span></td>
      </tr>
      <tr>
        <td id="L140" class="blob-num js-line-number" data-line-number="140"></td>
        <td id="LC140" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L141" class="blob-num js-line-number" data-line-number="141"></td>
        <td id="LC141" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L142" class="blob-num js-line-number" data-line-number="142"></td>
        <td id="LC142" class="blob-code blob-code-inner js-file-line"><span class="pl-c"><span class="pl-c">--</span> commands for bus unit</span></td>
      </tr>
      <tr>
        <td id="L143" class="blob-num js-line-number" data-line-number="143"></td>
        <td id="LC143" class="blob-code blob-code-inner js-file-line"><span class="pl-k">type</span> <span class="pl-en">busops_t</span> <span class="pl-k">is</span> (BUS_READB, BUS_READBU, BUS_READH, BUS_READHU, BUS_READW, BUS_WRITEB, BUS_WRITEH, BUS_WRITEW);</td>
      </tr>
      <tr>
        <td id="L144" class="blob-num js-line-number" data-line-number="144"></td>
        <td id="LC144" class="blob-code blob-code-inner js-file-line"><span class="pl-k">attribute</span> enum_encoding <span class="pl-k">of</span> busops_t : <span class="pl-k">type</span> <span class="pl-k">is</span> <span class="pl-s"><span class="pl-pds">&quot;</span>one-hot<span class="pl-pds">&quot;</span></span>;</td>
      </tr>
      <tr>
        <td id="L145" class="blob-num js-line-number" data-line-number="145"></td>
        <td id="LC145" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L146" class="blob-num js-line-number" data-line-number="146"></td>
        <td id="LC146" class="blob-code blob-code-inner js-file-line"><span class="pl-c"><span class="pl-c">--</span> commands for program counter unit (PCU)</span></td>
      </tr>
      <tr>
        <td id="L147" class="blob-num js-line-number" data-line-number="147"></td>
        <td id="LC147" class="blob-code blob-code-inner js-file-line"><span class="pl-k">type</span> <span class="pl-en">pcuops_t</span> <span class="pl-k">is</span> (PCU_SETPC, PCU_ENTERTRAP, PCU_RETTRAP, PCU_ENTERINT, PCU_RETINT);</td>
      </tr>
      <tr>
        <td id="L148" class="blob-num js-line-number" data-line-number="148"></td>
        <td id="LC148" class="blob-code blob-code-inner js-file-line"><span class="pl-k">attribute</span> enum_encoding <span class="pl-k">of</span> pcuops_t : <span class="pl-k">type</span> <span class="pl-k">is</span> <span class="pl-s"><span class="pl-pds">&quot;</span>one-hot<span class="pl-pds">&quot;</span></span>;</td>
      </tr>
      <tr>
        <td id="L149" class="blob-num js-line-number" data-line-number="149"></td>
        <td id="LC149" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L150" class="blob-num js-line-number" data-line-number="150"></td>
        <td id="LC150" class="blob-code blob-code-inner js-file-line"><span class="pl-c"><span class="pl-c">--</span> commands for register unit</span></td>
      </tr>
      <tr>
        <td id="L151" class="blob-num js-line-number" data-line-number="151"></td>
        <td id="LC151" class="blob-code blob-code-inner js-file-line"><span class="pl-k">type</span> <span class="pl-en">regops_t</span> <span class="pl-k">is</span> (REGOP_READ, REGOP_WRITE);</td>
      </tr>
      <tr>
        <td id="L152" class="blob-num js-line-number" data-line-number="152"></td>
        <td id="LC152" class="blob-code blob-code-inner js-file-line"><span class="pl-k">attribute</span> enum_encoding <span class="pl-k">of</span> regops_t : <span class="pl-k">type</span> <span class="pl-k">is</span> <span class="pl-s"><span class="pl-pds">&quot;</span>sequential<span class="pl-pds">&quot;</span></span>;</td>
      </tr>
      <tr>
        <td id="L153" class="blob-num js-line-number" data-line-number="153"></td>
        <td id="LC153" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L154" class="blob-num js-line-number" data-line-number="154"></td>
        <td id="LC154" class="blob-code blob-code-inner js-file-line"><span class="pl-k">end</span> <span class="pl-en">constants</span>;</td>
      </tr>
      <tr>
        <td id="L155" class="blob-num js-line-number" data-line-number="155"></td>
        <td id="LC155" class="blob-code blob-code-inner js-file-line">
</td>
      </tr>
      <tr>
        <td id="L156" class="blob-num js-line-number" data-line-number="156"></td>
        <td id="LC156" class="blob-code blob-code-inner js-file-line"><span class="pl-k">package</span> <span class="pl-k">body</span> <span class="pl-en">constants</span> <span class="pl-k">is</span></td>
      </tr>
      <tr>
        <td id="L157" class="blob-num js-line-number" data-line-number="157"></td>
        <td id="LC157" class="blob-code blob-code-inner js-file-line"> </td>
      </tr>
      <tr>
        <td id="L158" class="blob-num js-line-number" data-line-number="158"></td>
        <td id="LC158" class="blob-code blob-code-inner js-file-line"><span class="pl-k">end</span> <span class="pl-en">constants</span>;</td>
      </tr>
</table>

  </div>

</div>

<button type="button" data-facebox="#jump-to-line" data-facebox-class="linejump" data-hotkey="l" class="d-none">Jump to Line</button>
<div id="jump-to-line" style="display:none">
  <!-- '"` --><!-- </textarea></xmp> --></option></form><form accept-charset="UTF-8" action="" class="js-jump-to-line-form" method="get"><div style="margin:0;padding:0;display:inline"><input name="utf8" type="hidden" value="&#x2713;" /></div>
    <input class="form-control linejump-input js-jump-to-line-field" type="text" placeholder="Jump to line&hellip;" aria-label="Jump to line" autofocus>
    <button type="submit" class="btn">Go</button>
</form></div>


  </div>
  <div class="modal-backdrop js-touch-events"></div>
</div>

    </div>
  </div>

  </div>

      
<div class="container site-footer-container">
  <div class="site-footer " role="contentinfo">
    <ul class="site-footer-links float-right">
        <li><a href="https://github.com/contact" data-ga-click="Footer, go to contact, text:contact">Contact GitHub</a></li>
      <li><a href="https://developer.github.com" data-ga-click="Footer, go to api, text:api">API</a></li>
      <li><a href="https://training.github.com" data-ga-click="Footer, go to training, text:training">Training</a></li>
      <li><a href="https://shop.github.com" data-ga-click="Footer, go to shop, text:shop">Shop</a></li>
        <li><a href="https://github.com/blog" data-ga-click="Footer, go to blog, text:blog">Blog</a></li>
        <li><a href="https://github.com/about" data-ga-click="Footer, go to about, text:about">About</a></li>

    </ul>

    <a href="https://github.com" aria-label="Homepage" class="site-footer-mark" title="GitHub">
      <svg aria-hidden="true" class="octicon octicon-mark-github" height="24" version="1.1" viewBox="0 0 16 16" width="24"><path fill-rule="evenodd" d="M8 0C3.58 0 0 3.58 0 8c0 3.54 2.29 6.53 5.47 7.59.4.07.55-.17.55-.38 0-.19-.01-.82-.01-1.49-2.01.37-2.53-.49-2.69-.94-.09-.23-.48-.94-.82-1.13-.28-.15-.68-.52-.01-.53.63-.01 1.08.58 1.23.82.72 1.21 1.87.87 2.33.66.07-.52.28-.87.51-1.07-1.78-.2-3.64-.89-3.64-3.95 0-.87.31-1.59.82-2.15-.08-.2-.36-1.02.08-2.12 0 0 .67-.21 2.2.82.64-.18 1.32-.27 2-.27.68 0 1.36.09 2 .27 1.53-1.04 2.2-.82 2.2-.82.44 1.1.16 1.92.08 2.12.51.56.82 1.27.82 2.15 0 3.07-1.87 3.75-3.65 3.95.29.25.54.73.54 1.48 0 1.07-.01 1.93-.01 2.2 0 .21.15.46.55.38A8.013 8.013 0 0 0 16 8c0-4.42-3.58-8-8-8z"/></svg>
</a>
    <ul class="site-footer-links">
      <li>&copy; 2017 <span title="0.13137s from github-fe151-cp1-prd.iad.github.net">GitHub</span>, Inc.</li>
        <li><a href="https://github.com/site/terms" data-ga-click="Footer, go to terms, text:terms">Terms</a></li>
        <li><a href="https://github.com/site/privacy" data-ga-click="Footer, go to privacy, text:privacy">Privacy</a></li>
        <li><a href="https://github.com/security" data-ga-click="Footer, go to security, text:security">Security</a></li>
        <li><a href="https://status.github.com/" data-ga-click="Footer, go to status, text:status">Status</a></li>
        <li><a href="https://help.github.com" data-ga-click="Footer, go to help, text:help">Help</a></li>
    </ul>
  </div>
</div>



  

  <div id="ajax-error-message" class="ajax-error-message flash flash-error">
    <svg aria-hidden="true" class="octicon octicon-alert" height="16" version="1.1" viewBox="0 0 16 16" width="16"><path fill-rule="evenodd" d="M8.865 1.52c-.18-.31-.51-.5-.87-.5s-.69.19-.87.5L.275 13.5c-.18.31-.18.69 0 1 .19.31.52.5.87.5h13.7c.36 0 .69-.19.86-.5.17-.31.18-.69.01-1L8.865 1.52zM8.995 13h-2v-2h2v2zm0-3h-2V6h2v4z"/></svg>
    <button type="button" class="flash-close js-flash-close js-ajax-error-dismiss" aria-label="Dismiss error">
      <svg aria-hidden="true" class="octicon octicon-x" height="16" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M7.48 8l3.75 3.75-1.48 1.48L6 9.48l-3.75 3.75-1.48-1.48L4.52 8 .77 4.25l1.48-1.48L6 6.52l3.75-3.75 1.48 1.48z"/></svg>
    </button>
    You can't perform that action at this time.
  </div>


    
    <script crossorigin="anonymous" integrity="sha256-X+Q/xqnlEgxCczSjjpp2AUGGgqM5gcBzhRQ0p+EAUEk=" src="https://assets-cdn.github.com/assets/frameworks-5fe43fc6a9e5120c427334a38e9a7601418682a33981c073851434a7e1005049.js"></script>
    <script async="async" crossorigin="anonymous" integrity="sha256-9juSBU/6LfdytN4FT9IaLZ+xufYSqHkBZRUgHcrSaCw=" src="https://assets-cdn.github.com/assets/github-f63b92054ffa2df772b4de054fd21a2d9fb1b9f612a879016515201dcad2682c.js"></script>
    
    
    
    
  <div class="js-stale-session-flash stale-session-flash flash flash-warn flash-banner d-none">
    <svg aria-hidden="true" class="octicon octicon-alert" height="16" version="1.1" viewBox="0 0 16 16" width="16"><path fill-rule="evenodd" d="M8.865 1.52c-.18-.31-.51-.5-.87-.5s-.69.19-.87.5L.275 13.5c-.18.31-.18.69 0 1 .19.31.52.5.87.5h13.7c.36 0 .69-.19.86-.5.17-.31.18-.69.01-1L8.865 1.52zM8.995 13h-2v-2h2v2zm0-3h-2V6h2v4z"/></svg>
    <span class="signed-in-tab-flash">You signed in with another tab or window. <a href="">Reload</a> to refresh your session.</span>
    <span class="signed-out-tab-flash">You signed out in another tab or window. <a href="">Reload</a> to refresh your session.</span>
  </div>
  <div class="facebox" id="facebox" style="display:none;">
  <div class="facebox-popup">
    <div class="facebox-content" role="dialog" aria-labelledby="facebox-header" aria-describedby="facebox-description">
    </div>
    <button type="button" class="facebox-close js-facebox-close" aria-label="Close modal">
      <svg aria-hidden="true" class="octicon octicon-x" height="16" version="1.1" viewBox="0 0 12 16" width="12"><path fill-rule="evenodd" d="M7.48 8l3.75 3.75-1.48 1.48L6 9.48l-3.75 3.75-1.48-1.48L4.52 8 .77 4.25l1.48-1.48L6 6.52l3.75-3.75 1.48 1.48z"/></svg>
    </button>
  </div>
</div>


  </body>
</html>

